-- Elementos de Sistemas
-- by Luciano Soares
-- ALU.vhd

-- Unidade Lógica Aritmética (ULA)
-- Recebe dois valores de 16bits e
-- calcula uma das seguintes funções:
-- X+y, x-y, y-x, 0, 1, -1, x, y, -x, -y,
-- X+1, y+1, x-1, y-1, x&y, x|y
-- De acordo com os 6 bits de entrada denotados:
-- zx, nx, zy, ny, f, no.
-- Também calcula duas saídas de 1 bit:
-- Se a saída == 0, zr é definida como 1, senão 0;
-- Se a saída <0, ng é definida como 1, senão 0.
-- a ULA opera sobre os valores, da seguinte forma:
-- se (zx == 1) então x = 0
-- se (nx == 1) então x =! X
-- se (zy == 1) então y = 0
-- se (ny == 1) então y =! Y
-- se (f == 1) então saída = x + y
-- se (f == 0) então saída = x & y
-- se (no == 1) então saída = !saída
-- se (out == 0) então zr = 1
-- se (out <0) então ng = 1

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ALU is
	port (
			x,y:   in STD_LOGIC_VECTOR(15 downto 0); -- entradas de dados da ALU
			zx:    in STD_LOGIC;                     -- zera a entrada x
			nx:    in STD_LOGIC;                     -- inverte a entrada x
			zy:    in STD_LOGIC;                     -- zera a entrada y
			ny:    in STD_LOGIC;                     -- inverte a entrada y
			f:     in STD_LOGIC_VECTOR(1 downto 0);  -- se 0 calcula x & y, senão x + y
			no:    in STD_LOGIC;                     -- inverte o valor da saída
			zr:    out STD_LOGIC;                    -- setado se saída igual a zero
			ng:    out STD_LOGIC;                    -- setado se saída é negativa
			saida: out STD_LOGIC_VECTOR(15 downto 0) -- saída de dados da ALU
	);
end entity;

architecture  rtl OF alu is
  -- Aqui declaramos sinais (fios auxiliares)
  -- e componentes (outros módulos) que serao
  -- utilizados nesse modulo.

	component zerador16 IS
		port(z   : in STD_LOGIC;
			 a   : in STD_LOGIC_VECTOR(15 downto 0);
			 y   : out STD_LOGIC_VECTOR(15 downto 0)
			);
	end component;

	component inversor16 is
		port(z   : in STD_LOGIC;
			 a   : in STD_LOGIC_VECTOR(15 downto 0);
			 y   : out STD_LOGIC_VECTOR(15 downto 0)
		);
	end component;

	component Add16 is
		port(
			a   :  in STD_LOGIC_VECTOR(15 downto 0);
			b   :  in STD_LOGIC_VECTOR(15 downto 0);
			q   : out STD_LOGIC_VECTOR(15 downto 0)
		);
	end component;

	component BarrelShifter16 is
		port ( 
			a:    in  STD_LOGIC_VECTOR(15 downto 0);   -- input vector
			dir:  in  STD_LOGIC;                       -- 0=>left 1=>right
			size: in  STD_LOGIC_VECTOR(2 downto 0);    -- shift amount
			q:    out STD_LOGIC_VECTOR(15 downto 0)    -- output vector (shifted)
		);
	end component;

	component comparador16 is
		port(
			a    : in STD_LOGIC_VECTOR(15 downto 0);
			zr   : out STD_LOGIC;                  
			ng   : out STD_LOGIC
   		 );
	end component;

	component Mux4Way16 is
		port (
			a:   in  STD_LOGIC_VECTOR(15 downto 0);
			b:   in  STD_LOGIC_VECTOR(15 downto 0);
			c:   in  STD_LOGIC_VECTOR(15 downto 0);
			D:   in  STD_LOGIC_VECTOR(15 downto 0);
			sel: in  STD_LOGIC_VECTOR(1 downto 0);
			q:   out STD_LOGIC_VECTOR(15 downto 0)
		);
	end component;
	
   SIGNAL zxout,zyout,nxout,nyout,andout,adderout,barrelout,muxout,precomp: std_logic_vector(15 downto 0);	

--    when zx = '0' zxout <= x else zxout <= "0000000000000000";
--    when nx = '0' nxout <= zxout else nxout <= !zxout;
--    when zy = '0' zyout <= y else zyout <= "0000000000000000";
--    when ny = '0' nyout <= zyout else nyout <= !zyout;
--    andout <= nxout and nyout;
--    adderout <= 
begin
    -- Implementação vem aqui!
	z1: zerador16 port map (
		z => zx,
		a => x,
		y => zxout
	);

	z2: zerador16 port map (
		z => zy,
		a => y,
		y => zyout
	);

	i1: inversor16 port map (	
		z => nx,
		a => zxout,
		y => nxout
	);

	i2: inversor16 port map (	
		z => ny,
		a => zyout,
		y => nyout
	);

	andout <= nxout and nyout;

	add: Add16 port map (
		a => nxout,
		b => nyout,
		q => adderout
	);

	multiplica: BarrelShifter16 port map(
		a => nxout,
		dir => f(0),
		size => "001",
		q => barrelout
	);

	mux: Mux4Way16 port map(
		a => andout,
		b => adderout,
		c => barrelout,
		d => barrelout,
		sel => f,
		q => muxout
	);

	i3: inversor16 port map (	
		z => no,
		a => muxout,
		y => precomp
	);

	saida <= precomp;

	comp: comparador16 port map (
		a => precomp,                                                      
		zr => zr,
		ng => ng
	);

end architecture;
